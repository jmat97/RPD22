/**
 * Copyright (C) 2020  AGH University of Science and Technology
 *
 * This program is free software: you can redistribute it and/or modify
 * it under the terms of the GNU General Public License as published by
 * the Free Software Foundation, either version 3 of the License, or
 * (at your option) any later version.
 *
 * This program is distributed in the hope that it will be useful,
 * but WITHOUT ANY WARRANTY; without even the implied warranty of
 * MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
 * GNU General Public License for more details.
 *
 * You should have received a copy of the GNU General Public License
 * along with this program.  If not, see <https://www.gnu.org/licenses/>.
 */

interface rst_if (
    output logic rst_n,
    input logic  clk
);


/**
 * Tasks and functions definitions
 */

function void init();
    rst_n = 1'b1;
endfunction

task reset();
    @(posedge clk) ;
    @(negedge clk) ;
    rst_n = 1'b0;
    @(negedge clk) ;
    rst_n = 1'b1;
endtask

endinterface
